DATE,EXERCISE,NB_REPS,WEIGHT,DURATION
06-06-2022,Extensions triceps 1 haltère,12,20.0,00:00:00
06-06-2022,Curl concentré,12,20.0,00:00:00
06-06-2022,Extensions triceps 1 haltère,15,18.0,00:00:00
06-06-2022,Curl barre,12,40.0,00:00:00
06-06-2022,Curl barre,12,40.0,00:00:00
06-06-2022,Curl barre,12,40.0,00:00:00
06-06-2022,Curl barre,15,30.0,00:00:00
30-05-2022,Gainage,0,PDC,00:01:30
30-05-2022,Gainage,0,PDC,00:02:30
30-05-2022,Gainage,0,PDC,00:02:30
30-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
30-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
30-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
30-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
30-05-2022,[Basic] Seated dip,12,77.0,00:00:00
30-05-2022,[Basic] Seated dip,12,77.0,00:00:00
30-05-2022,[Basic] Seated dip,12,77.0,00:00:00
30-05-2022,[Basic] Seated dip,12,77.0,00:00:00
30-05-2022,[Basic] Arm curl,11,54.0,00:00:00
30-05-2022,[Basic] Arm curl,11,54.0,00:00:00
30-05-2022,[Basic] Arm curl,11,54.0,00:00:00
30-05-2022,[Basic] Arm curl,11,54.0,00:00:00
30-05-2022,Curl concentré,11,20.0,00:00:00
30-05-2022,Extensions triceps 1 haltère,11,20.0,00:00:00
30-05-2022,Extensions triceps 1 haltère,11,20.0,00:00:00
30-05-2022,Extensions triceps 1 haltère,11,20.0,00:00:00
30-05-2022,Extensions triceps 1 haltère,11,20.0,00:00:00
30-05-2022,Curl concentré,11,20.0,00:00:00
30-05-2022,Curl concentré,11,20.0,00:00:00
30-05-2022,Curl concentré,11,20.0,00:00:00
30-05-2022,Barre au front derriere la tête,11,32.0,00:00:00
30-05-2022,Curl barre,11,40.0,00:00:00
30-05-2022,Curl barre,11,40.0,00:00:00
30-05-2022,Barre au front derriere la tête,11,32.0,00:00:00
30-05-2022,Barre au front derriere la tête,12,30.0,00:00:00
30-05-2022,Barre au front derriere la tête,12,30.0,00:00:00
30-05-2022,Curl barre,11,40.0,00:00:00
30-05-2022,Curl barre,15,30.0,00:00:00
28-05-2022,[Basic] Abdominal,9,41.0,00:00:00
28-05-2022,[Basic] Abdominal,9,41.0,00:00:00
28-05-2022,[Basic] Abdominal,10,45.0,00:00:00
28-05-2022,[Basic] Abdominal,8,45.0,00:00:00
28-05-2022,Gainage,0,PDC,00:01:30
28-05-2022,Gainage,0,PDC,00:02:30
28-05-2022,Gainage,0,PDC,00:02:30
28-05-2022,[Basic] Lat pulldown,10,52.0,00:00:00
28-05-2022,[Basic] Lat pulldown,11,52.0,00:00:00
28-05-2022,[Basic] Lat pulldown,12,52.0,00:00:00
28-05-2022,[Basic] Lat pulldown,12,52.0,00:00:00
28-05-2022,[Basic] Diverging lat pulldown,8,52.0,00:00:00
28-05-2022,[Basic] Diverging lat pulldown,8,52.0,00:00:00
28-05-2022,[Basic] Diverging lat pulldown,8,52.0,00:00:00
28-05-2022,[Basic] Diverging lat pulldown,8,52.0,00:00:00
28-05-2022,Tirage menton haltères ,11,16.0,00:00:00
28-05-2022,Tirage menton haltères ,11,16.0,00:00:00
28-05-2022,Tirage menton haltères ,11,16.0,00:00:00
28-05-2022,Tirage menton haltères ,11,16.0,00:00:00
28-05-2022,Rowing barre,8,70.0,00:00:00
28-05-2022,Rowing barre,8,70.0,00:00:00
28-05-2022,Rowing barre,8,70.0,00:00:00
28-05-2022,Rowing barre,15,30.0,00:00:00
26-05-2022,Développé épaules à la machine,11,50.0,00:00:00
26-05-2022,Gainage,0,PDC,00:01:30
26-05-2022,Gainage,0,PDC,00:02:30
26-05-2022,Gainage,0,PDC,00:02:30
26-05-2022,[Basic] Abdominal crunch,12,82.0,00:00:00
26-05-2022,[Basic] Abdominal crunch,12,82.0,00:00:00
26-05-2022,[Basic] Abdominal crunch,12,82.0,00:00:00
26-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
26-05-2022,Élévations latérales,10,9.0,00:00:00
26-05-2022,Élévations latérales,10,9.0,00:00:00
26-05-2022,Élévations latérales,10,9.0,00:00:00
26-05-2022,Élévations latérales,10,9.0,00:00:00
26-05-2022,Développé Arnold,10,16.0,00:00:00
26-05-2022,Développé Arnold,10,16.0,00:00:00
26-05-2022,Développé Arnold,10,16.0,00:00:00
26-05-2022,Développé Arnold,10,16.0,00:00:00
26-05-2022,Développé militaire haltères,8,24.0,00:00:00
26-05-2022,Développé militaire haltères,8,24.0,00:00:00
26-05-2022,Développé militaire haltères,11,24.0,00:00:00
26-05-2022,Développé militaire haltères,11,24.0,00:00:00
26-05-2022,Développé militaire haltères,20,16.0,00:00:00
24-05-2022,[Basic] Chest press,8,59.0,00:00:00
24-05-2022,[Basic] Chest press,8,59.0,00:00:00
24-05-2022,[Basic] Chest press,8,59.0,00:00:00
24-05-2022,[Basic] Chest press,8,59.0,00:00:00
24-05-2022,Écarté Haltères,12,14.0,00:00:00
24-05-2022,Écarté Haltères,12,14.0,00:00:00
24-05-2022,Écarté Haltères,12,14.0,00:00:00
24-05-2022,Écarté Haltères,12,14.0,00:00:00
24-05-2022,Développé incliné,8,57.0,00:00:00
24-05-2022,Développé incliné,8,57.0,00:00:00
24-05-2022,Développé incliné,8,57.0,00:00:00
24-05-2022,Développé incliné,8,57.0,00:00:00
24-05-2022,Développé couché,10,60.0,00:00:00
24-05-2022,Développé couché,10,60.0,00:00:00
24-05-2022,Développé couché,10,60.0,00:00:00
24-05-2022,Développé couché,15,40.0,00:00:00
23-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
23-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
23-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
23-05-2022,[Basic] Arm curl,8,54.0,00:00:00
23-05-2022,[Basic] Seated dip,8,77.0,00:00:00
23-05-2022,[Basic] Seated dip,8,77.0,00:00:00
23-05-2022,[Basic] Arm curl,8,54.0,00:00:00
23-05-2022,[Basic] Arm curl,8,54.0,00:00:00
23-05-2022,[Basic] Seated dip,8,77.0,00:00:00
23-05-2022,[Basic] Seated dip,12,77.0,00:00:00
23-05-2022,[Basic] Arm curl,10,54.0,00:00:00
23-05-2022,Extensions triceps 1 haltère,11,18.0,00:00:00
23-05-2022,Extensions triceps 1 haltère,10,20.0,00:00:00
23-05-2022,Curl concentré,8,20.0,00:00:00
23-05-2022,Curl concentré,9,20.0,00:00:00
23-05-2022,Curl concentré,10,20.0,00:00:00
23-05-2022,Curl concentré,10,20.0,00:00:00
23-05-2022,Extensions triceps 1 haltère,10,20.0,00:00:00
23-05-2022,Extensions triceps 1 haltère,10,20.0,00:00:00
23-05-2022,Curl concentré,10,20.0,00:00:00
23-05-2022,Barre au front derriere la tête,10,32.0,00:00:00
23-05-2022,Curl barre,9,40.0,00:00:00
23-05-2022,Barre au front derriere la tête,7,35.0,00:00:00
23-05-2022,Barre au front derriere la tête,8,35.0,00:00:00
23-05-2022,Barre au front derriere la tête,15,30.0,00:00:00
23-05-2022,Curl barre,10,40.0,00:00:00
23-05-2022,Curl barre,10,40.0,00:00:00
23-05-2022,Curl barre,15,30.0,00:00:00
21-05-2022,Gainage,0,PDC,00:01:30
21-05-2022,Gainage,0,PDC,00:02:30
21-05-2022,Gainage,0,PDC,00:02:30
21-05-2022,[Basic] Abdominal crunch,6,82.0,00:00:00
21-05-2022,[Basic] Abdominal crunch,9,82.0,00:00:00
21-05-2022,[Basic] Abdominal crunch,9,82.0,00:00:00
21-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
21-05-2022,[Basic] Seated row,10,59.0,00:00:00
21-05-2022,[Basic] Seated row,10,59.0,00:00:00
21-05-2022,[Basic] Seated row,10,59.0,00:00:00
21-05-2022,[Basic] Seated row,10,59.0,00:00:00
21-05-2022,[Basic] Diverging lat pulldown,12,45.0,00:00:00
21-05-2022,[Basic] Diverging lat pulldown,12,45.0,00:00:00
21-05-2022,[Basic] Diverging lat pulldown,12,45.0,00:00:00
21-05-2022,[Basic] Diverging lat pulldown,12,45.0,00:00:00
21-05-2022,Tirage menton haltères ,10,16.0,00:00:00
21-05-2022,Tirage menton haltères ,10,16.0,00:00:00
21-05-2022,Tirage menton haltères ,10,16.0,00:00:00
21-05-2022,Tirage menton haltères ,10,16.0,00:00:00
21-05-2022,Rowing barre,8,70.0,00:00:00
21-05-2022,Rowing barre,12,60.0,00:00:00
21-05-2022,Rowing barre,12,50.0,00:00:00
21-05-2022,Rowing barre,15,30.0,00:00:00
19-05-2022,[Basic] Abdominal crunch,12,77.0,00:00:00
19-05-2022,[Basic] Abdominal crunch,12,77.0,00:00:00
19-05-2022,[Basic] Abdominal crunch,12,77.0,00:00:00
19-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
19-05-2022,Développé épaules à la machine,10,50.0,00:00:00
19-05-2022,Développé épaules à la machine,10,50.0,00:00:00
19-05-2022,Développé épaules à la machine,10,50.0,00:00:00
19-05-2022,Développé épaules à la machine,10,50.0,00:00:00
19-05-2022,Élévations latérales,9,9.0,00:00:00
19-05-2022,Élévations latérales,9,9.0,00:00:00
19-05-2022,Élévations latérales,9,9.0,00:00:00
19-05-2022,Élévations latérales,9,9.0,00:00:00
19-05-2022,Développé Arnold,9,16.0,00:00:00
19-05-2022,Développé Arnold,9,16.0,00:00:00
19-05-2022,Développé Arnold,9,16.0,00:00:00
19-05-2022,Développé Arnold,9,16.0,00:00:00
19-05-2022,Développé militaire haltères,10,22.0,00:00:00
19-05-2022,Développé militaire haltères,12,22.0,00:00:00
19-05-2022,Développé militaire haltères,12,22.0,00:00:00
19-05-2022,Développé militaire haltères,12,22.0,00:00:00
19-05-2022,Développé militaire haltères,15,14.0,00:00:00
17-05-2022,[Basic] Chest press,8,52.0,00:00:00
17-05-2022,[Basic] Chest press,8,52.0,00:00:00
17-05-2022,[Basic] Chest press,8,52.0,00:00:00
17-05-2022,[Basic] Chest press,8,55.0,00:00:00
17-05-2022,Butterfly,8,73.0,00:00:00
17-05-2022,Butterfly,8,73.0,00:00:00
17-05-2022,Butterfly,8,79.0,00:00:00
17-05-2022,Butterfly,9,79.0,00:00:00
17-05-2022,Écarté Haltères,11,14.0,00:00:00
17-05-2022,Écarté Haltères,11,14.0,00:00:00
17-05-2022,Écarté Haltères,11,14.0,00:00:00
17-05-2022,Écarté Haltères,11,14.0,00:00:00
17-05-2022,Développé couché,8,60.0,00:00:00
17-05-2022,Développé couché,8,60.0,00:00:00
17-05-2022,Développé couché,9,60.0,00:00:00
17-05-2022,Développé couché,9,60.0,00:00:00
17-05-2022,Développé incliné,9,55.0,00:00:00
17-05-2022,Développé incliné,9,55.0,00:00:00
17-05-2022,Développé incliné,9,55.0,00:00:00
17-05-2022,Développé incliné,16,40.0,00:00:00
16-05-2022,[Basic] Seated dip,12,73.0,00:00:00
16-05-2022,[Basic] Seated dip,12,73.0,00:00:00
16-05-2022,[Basic] Seated dip,12,73.0,00:00:00
16-05-2022,Curl supination barre,8,35.0,00:00:00
16-05-2022,Curl supination barre,8,35.0,00:00:00
16-05-2022,Curl supination barre,8,35.0,00:00:00
16-05-2022,Curl supination barre,12,30.0,00:00:00
16-05-2022,Extensions triceps 1 haltère,9,20.0,00:00:00
16-05-2022,Curl concentré,9,20.0,00:00:00
16-05-2022,Curl concentré,9,20.0,00:00:00
16-05-2022,Extensions triceps 1 haltère,9,20.0,00:00:00
16-05-2022,Extensions triceps 1 haltère,9,20.0,00:00:00
16-05-2022,Curl concentré,9,20.0,00:00:00
16-05-2022,Extensions triceps 1 haltère,12,18.0,00:00:00
16-05-2022,Curl concentré,9,20.0,00:00:00
16-05-2022,Barre au front derriere la tête,4,40.0,00:00:00
16-05-2022,Barre au front derriere la tête,12,30.0,00:00:00
16-05-2022,Barre au front derriere la tête,12,30.0,00:00:00
16-05-2022,Barre au front derriere la tête,15,25.0,00:00:00
16-05-2022,Curl barre,8,40.0,00:00:00
16-05-2022,Curl barre,9,40.0,00:00:00
16-05-2022,Curl barre,9,40.0,00:00:00
16-05-2022,Curl barre,12,30.0,00:00:00
14-05-2022,Gainage,0,PDC,00:01:30
14-05-2022,Gainage,0,PDC,00:02:30
14-05-2022,Gainage,0,PDC,00:02:30
14-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
14-05-2022,[Basic] Abdominal crunch,8,82.0,00:00:00
14-05-2022,[Basic] Abdominal crunch,8,82.0,00:00:00
14-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
14-05-2022,Tractions nuque,8,PDC,00:00:00
14-05-2022,Tractions nuque,8,PDC,00:00:00
14-05-2022,Tractions nuque,8,PDC,00:00:00
14-05-2022,Tractions nuque,8,PDC,00:00:00
14-05-2022,[Basic] Lat pulldown,11,52.0,00:00:00
14-05-2022,[Basic] Lat pulldown,11,52.0,00:00:00
14-05-2022,[Basic] Lat pulldown,11,52.0,00:00:00
14-05-2022,[Basic] Lat pulldown,11,52.0,00:00:00
14-05-2022,Tirage menton haltères ,9,16.0,00:00:00
14-05-2022,Tirage menton haltères ,9,16.0,00:00:00
14-05-2022,Tirage menton haltères ,9,16.0,00:00:00
14-05-2022,Tirage menton haltères ,9,16.0,00:00:00
14-05-2022,Rowing barre,12,50.0,00:00:00
14-05-2022,Rowing barre,12,50.0,00:00:00
14-05-2022,Rowing barre,12,50.0,00:00:00
14-05-2022,Rowing barre,15,30.0,00:00:00
10-05-2022,Gainage,0,PDC,00:01:15
10-05-2022,Gainage,0,PDC,00:02:15
10-05-2022,Gainage,0,PDC,00:02:15
10-05-2022,[Basic] Abdominal crunch,12,68.0,00:00:00
10-05-2022,[Basic] Abdominal crunch,12,77.0,00:00:00
10-05-2022,[Basic] Abdominal crunch,12,77.0,00:00:00
10-05-2022,[Basic] Abdominal crunch,10,73.0,00:00:00
10-05-2022,Butterfly,8,73.0,00:00:00
10-05-2022,Butterfly,8,73.0,00:00:00
10-05-2022,Butterfly,8,79.0,00:00:00
10-05-2022,Butterfly,9,79.0,00:00:00
10-05-2022,[Basic] Chest press,8,59.0,00:00:00
10-05-2022,[Basic] Chest press,8,59.0,00:00:00
10-05-2022,[Basic] Chest press,8,59.0,00:00:00
10-05-2022,[Basic] Chest press,9,59.0,00:00:00
10-05-2022,Écarté Haltères,10,14.0,00:00:00
10-05-2022,Écarté Haltères,10,14.0,00:00:00
10-05-2022,Écarté Haltères,10,14.0,00:00:00
10-05-2022,Écarté Haltères,10,14.0,00:00:00
10-05-2022,Développé couché avec haltères,9,22.0,00:00:00
10-05-2022,Développé couché avec haltères,9,22.0,00:00:00
10-05-2022,Développé couché avec haltères,11,22.0,00:00:00
10-05-2022,Développé couché avec haltères,11,22.0,00:00:00
10-05-2022,Développé incliné,8,55.0,00:00:00
10-05-2022,Développé incliné,8,55.0,00:00:00
10-05-2022,Développé incliné,8,55.0,00:00:00
10-05-2022,Développé incliné,12,50.0,00:00:00
10-05-2022,Développé incliné,17,20.0,00:00:00
09-05-2022,[Basic] Seated dip,12,68.0,00:00:00
09-05-2022,[Basic] Seated dip,12,68.0,00:00:00
09-05-2022,[Basic] Seated dip,12,68.0,00:00:00
09-05-2022,[Basic] Seated dip,10,68.0,00:00:00
09-05-2022,[Basic] Arm curl,12,50.0,00:00:00
09-05-2022,[Basic] Arm curl,12,50.0,00:00:00
09-05-2022,[Basic] Arm curl,12,50.0,00:00:00
09-05-2022,[Basic] Arm curl,12,45.0,00:00:00
09-05-2022,Dips,11,PDC,00:00:00
09-05-2022,Dips,15,PDC,00:00:00
09-05-2022,Dips,13,PDC,00:00:00
09-05-2022,Dips,15,PDC,00:00:00
09-05-2022,Curl supination barre,9,30.0,00:00:00
09-05-2022,Curl supination barre,12,30.0,00:00:00
09-05-2022,Curl supination barre,12,30.0,00:00:00
09-05-2022,Curl supination barre,12,30.0,00:00:00
09-05-2022,Extensions triceps 1 haltère,12,18.0,00:00:00
09-05-2022,Extensions triceps 1 haltère,12,18.0,00:00:00
09-05-2022,Extensions triceps 1 haltère,12,18.0,00:00:00
09-05-2022,Extensions triceps 1 haltère,12,18.0,00:00:00
09-05-2022,Curl barre,8,40.0,00:00:00
09-05-2022,Curl barre,8,40.0,00:00:00
09-05-2022,Curl barre,8,40.0,00:00:00
09-05-2022,Curl barre,12,30.0,00:00:00
07-05-2022,[Basic] Rameur,12,45.0,00:00:00
07-05-2022,[Basic] Rameur,12,45.0,00:00:00
07-05-2022,[Basic] Rameur,12,45.0,00:00:00
07-05-2022,[Basic] Rameur,12,45.0,00:00:00
07-05-2022,Gainage,0,PDC,00:01:15
07-05-2022,Gainage,0,PDC,00:02:15
07-05-2022,Gainage,0,PDC,00:02:15
07-05-2022,Tractions nuque,8,PDC,00:00:00
07-05-2022,Tractions nuque,8,PDC,00:00:00
07-05-2022,Tractions nuque,8,PDC,00:00:00
07-05-2022,Tractions nuque,9,PDC,00:00:00
07-05-2022,Tirage menton haltères ,8,16.0,00:00:00
07-05-2022,Tirage menton haltères ,8,16.0,00:00:00
07-05-2022,Tirage menton haltères ,8,16.0,00:00:00
07-05-2022,Tirage menton haltères ,8,16.0,00:00:00
07-05-2022,Rowing barre,11,60.0,00:00:00
07-05-2022,Rowing barre,11,60.0,00:00:00
07-05-2022,Rowing barre,11,60.0,00:00:00
07-05-2022,Rowing barre,12,30.0,00:00:00
05-05-2022,Développé épaules à la machine,9,50.0,00:00:00
05-05-2022,Développé épaules à la machine,9,50.0,00:00:00
05-05-2022,Développé épaules à la machine,9,50.0,00:00:00
05-05-2022,Gainage,0,PDC,00:01:15
05-05-2022,Gainage,0,PDC,00:02:15
05-05-2022,Gainage,0,PDC,00:02:15
05-05-2022,[Basic] Abdominal crunch,12,82.0,00:00:00
05-05-2022,[Basic] Abdominal crunch,11,82.0,00:00:00
05-05-2022,[Basic] Abdominal crunch,11,82.0,00:00:00
05-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
05-05-2022,Élévations latérales,9,9.0,00:00:00
05-05-2022,Élévations latérales,9,9.0,00:00:00
05-05-2022,Élévations latérales,9,9.0,00:00:00
05-05-2022,Élévations latérales,9,9.0,00:00:00
05-05-2022,Développé Arnold,8,16.0,00:00:00
05-05-2022,Développé Arnold,8,16.0,00:00:00
05-05-2022,Développé Arnold,8,16.0,00:00:00
05-05-2022,Développé Arnold,8,16.0,00:00:00
05-05-2022,Développé militaire haltères,12,22.0,00:00:00
05-05-2022,Développé militaire haltères,12,22.0,00:00:00
05-05-2022,Développé militaire haltères,12,22.0,00:00:00
05-05-2022,Développé militaire haltères,12,20.0,00:00:00
03-05-2022,Butterfly,7,79.0,00:00:00
03-05-2022,Butterfly,9,79.0,00:00:00
03-05-2022,[Basic] Converging chest press,7,52.0,00:00:00
03-05-2022,[Basic] Converging chest press,8,52.0,00:00:00
03-05-2022,[Basic] Converging chest press,8,52.0,00:00:00
03-05-2022,[Basic] Converging chest press,12,39.0,00:00:00
03-05-2022,Écarté Haltères,9,14.0,00:00:00
03-05-2022,Écarté Haltères,9,14.0,00:00:00
03-05-2022,Écarté Haltères,9,14.0,00:00:00
03-05-2022,Écarté Haltères,9,14.0,00:00:00
03-05-2022,Développé couché avec haltères,12,20.0,00:00:00
03-05-2022,Développé couché avec haltères,12,20.0,00:00:00
03-05-2022,Développé couché avec haltères,12,20.0,00:00:00
03-05-2022,Développé couché avec haltères,12,20.0,00:00:00
03-05-2022,Développé incliné avec haltères,12,20.0,00:00:00
03-05-2022,Développé couché,8,60.0,00:00:00
03-05-2022,Développé couché,9,60.0,00:00:00
03-05-2022,Développé couché,9,60.0,00:00:00
03-05-2022,Développé couché,15,40.0,00:00:00
02-05-2022,Gainage,0,PDC,00:01:15
02-05-2022,Gainage,0,PDC,00:02:15
02-05-2022,Gainage,0,PDC,00:02:15
02-05-2022,[Basic] Abdominal crunch,8,82.0,00:00:00
02-05-2022,[Basic] Abdominal crunch,8,82.0,00:00:00
02-05-2022,[Basic] Abdominal crunch,9,82.0,00:00:00
02-05-2022,[Basic] Abdominal crunch,12,73.0,00:00:00
02-05-2022,Curl biceps à la poulie basse,9,41.0,00:00:00
02-05-2022,Extension triceps poulie,8,45.0,00:00:00
02-05-2022,Extension triceps poulie,9,45.0,00:00:00
02-05-2022,Curl biceps à la poulie basse,10,41.0,00:00:00
02-05-2022,Curl biceps à la poulie basse,11,41.0,00:00:00
02-05-2022,Extension triceps poulie,9,45.0,00:00:00
02-05-2022,Extension triceps poulie,10,45.0,00:00:00
02-05-2022,Curl biceps à la poulie basse,11,41.0,00:00:00
02-05-2022,Extensions triceps 1 haltère,9,18.0,00:00:00
02-05-2022,Curl concentré,8,20.0,00:00:00
02-05-2022,Curl concentré,8,20.0,00:00:00
02-05-2022,Extensions triceps 1 haltère,9,18.0,00:00:00
02-05-2022,Extensions triceps 1 haltère,9,18.0,00:00:00
02-05-2022,Extensions triceps 1 haltère,10,18.0,00:00:00
02-05-2022,Curl concentré,8,20.0,00:00:00
02-05-2022,Curl concentré,9,20.0,00:00:00
02-05-2022,Barre au front derriere la tête,8,30.0,00:00:00
02-05-2022,Barre au front derriere la tête,8,30.0,00:00:00
02-05-2022,Barre au front derriere la tête,11,30.0,00:00:00
02-05-2022,Barre au front derriere la tête,12,30.0,00:00:00
02-05-2022,Curl barre,8,40.0,00:00:00
02-05-2022,Curl barre,8,40.0,00:00:00
02-05-2022,Curl barre,8,40.0,00:00:00
02-05-2022,Curl barre,12,30.0,00:00:00
30-04-2022,[Basic] Abdominal crunch,12,59.0,00:00:00
30-04-2022,[Basic] Abdominal crunch,12,72.0,00:00:00
30-04-2022,[Basic] Seated row,9,59.0,00:00:00
30-04-2022,[Basic] Seated row,9,59.0,00:00:00
30-04-2022,[Basic] Seated row,9,59.0,00:00:00
30-04-2022,[Basic] Seated row,9,59.0,00:00:00
30-04-2022,[Basic] Diverging lat pulldown,8,45.0,00:00:00
30-04-2022,[Basic] Diverging lat pulldown,8,45.0,00:00:00
30-04-2022,[Basic] Diverging lat pulldown,12,41.0,00:00:00
30-04-2022,[Basic] Diverging lat pulldown,12,41.0,00:00:00
30-04-2022,[Basic] Lat pulldown,10,52.0,00:00:00
30-04-2022,[Basic] Lat pulldown,10,52.0,00:00:00
30-04-2022,[Basic] Lat pulldown,10,52.0,00:00:00
30-04-2022,[Basic] Lat pulldown,10,52.0,00:00:00
30-04-2022,Tirage menton haltères ,12,14.0,00:00:00
30-04-2022,Tirage menton haltères ,12,14.0,00:00:00
30-04-2022,Tirage menton haltères ,12,14.0,00:00:00
30-04-2022,Tirage menton haltères ,12,14.0,00:00:00
30-04-2022,Rowing barre,10,60.0,00:00:00
30-04-2022,Rowing barre,10,60.0,00:00:00
30-04-2022,Rowing barre,10,60.0,00:00:00
30-04-2022,Rowing barre,12,30.0,00:00:00
28-04-2022,[Basic] Abdominal crunch,9,82.0,00:00:00
28-04-2022,[Basic] Abdominal crunch,12,77.0,00:00:00
28-04-2022,Gainage,0,PDC,00:01:00
28-04-2022,Gainage,0,PDC,00:01:30
28-04-2022,Gainage,0,PDC,00:02:00
28-04-2022,Développé épaules à la machine,6,50.0,00:00:00
28-04-2022,Développé épaules à la machine,8,50.0,00:00:00
28-04-2022,Développé épaules à la machine,8,50.0,00:00:00
28-04-2022,Développé épaules à la machine,8,50.0,00:00:00
28-04-2022,Élévations latérales,8,9.0,00:00:00
28-04-2022,Élévations latérales,8,9.0,00:00:00
28-04-2022,Élévations latérales,8,9.0,00:00:00
28-04-2022,Élévations latérales,8,9.0,00:00:00
28-04-2022,Développé Arnold,8,16.0,00:00:00
28-04-2022,Développé Arnold,8,16.0,00:00:00
28-04-2022,Développé Arnold,8,16.0,00:00:00
28-04-2022,Développé Arnold,8,16.0,00:00:00
28-04-2022,Développé militaire haltères,10,22.0,00:00:00
28-04-2022,Développé militaire haltères,10,22.0,00:00:00
28-04-2022,Développé militaire haltères,10,22.0,00:00:00
28-04-2022,Développé militaire haltères,12,20.0,00:00:00
26-04-2022,Gainage,0,PDC,00:01:30
26-04-2022,Gainage,0,PDC,00:02:00
26-04-2022,Gainage,0,PDC,00:02:00
26-04-2022,Développé épaules à la machine,8,41.0,00:00:00
26-04-2022,Développé épaules à la machine,8,41.0,00:00:00
26-04-2022,Développé épaules à la machine,7,45.0,00:00:00
26-04-2022,Développé épaules à la machine,7,50.0,00:00:00
26-04-2022,Butterfly,7,79.0,00:00:00
26-04-2022,Butterfly,8,79.0,00:00:00
26-04-2022,Butterfly,9,79.0,00:00:00
26-04-2022,Butterfly,12,73.0,00:00:00
26-04-2022,Élévations latérales,10,8.0,00:00:00
26-04-2022,Élévations latérales,10,8.0,00:00:00
26-04-2022,Élévations latérales,10,8.0,00:00:00
26-04-2022,Élévations latérales,8,8.0,00:00:00
26-04-2022,Écarté Haltères,8,14.0,00:00:00
26-04-2022,Développé militaire haltères,11,20.0,00:00:00
26-04-2022,Développé militaire haltères,11,20.0,00:00:00
26-04-2022,Écarté Haltères,8,14.0,00:00:00
26-04-2022,Écarté Haltères,8,14.0,00:00:00
26-04-2022,Développé incliné avec haltères,9,20.0,00:00:00
26-04-2022,Développé incliné avec haltères,9,20.0,00:00:00
26-04-2022,Développé incliné avec haltères,9,20.0,00:00:00
26-04-2022,Développé incliné avec haltères,9,20.0,00:00:00
26-04-2022,Développé couché avec haltères,8,22.0,00:00:00
26-04-2022,Développé couché avec haltères,9,22.0,00:00:00
26-04-2022,Développé couché avec haltères,12,22.0,00:00:00
26-04-2022,Développé couché avec haltères,12,20.0,00:00:00
25-04-2022,Gainage,0,PDC,00:01:00
25-04-2022,Gainage,0,PDC,00:02:00
25-04-2022,Gainage,0,PDC,00:02:00
25-04-2022,[Basic] Abdominal,10,41.0,00:00:00
25-04-2022,[Basic] Abdominal,10,41.0,00:00:00
25-04-2022,[Basic] Abdominal,10,41.0,00:00:00
25-04-2022,[Basic] Abdominal,10,41.0,00:00:00
25-04-2022,Extension triceps poulie,7,45.0,00:00:00
25-04-2022,Curl biceps à la poulie basse,8,41.0,00:00:00
25-04-2022,Extension triceps poulie,8,45.0,00:00:00
25-04-2022,Curl biceps à la poulie basse,8,41.0,00:00:00
25-04-2022,Extension triceps poulie,9,45.0,00:00:00
25-04-2022,Curl biceps à la poulie basse,12,36.0,00:00:00
25-04-2022,Extension triceps poulie,12,41.0,00:00:00
25-04-2022,Curl biceps à la poulie basse,12,32.0,00:00:00
25-04-2022,Extensions triceps 1 haltère,12,18.0,00:00:00
25-04-2022,Curl concentré,12,18.0,00:00:00
25-04-2022,Extensions triceps 1 haltère,12,18.0,00:00:00
25-04-2022,Curl concentré,12,18.0,00:00:00
25-04-2022,Extensions triceps 1 haltère,9,18.0,00:00:00
25-04-2022,Curl concentré,12,18.0,00:00:00
25-04-2022,Extensions triceps 1 haltère,9,18.0,00:00:00
25-04-2022,Curl concentré,12,18.0,00:00:00
25-04-2022,Barre au front derriere la tête,12,25.0,00:00:00
25-04-2022,Curl barre,12,30.0,00:00:00
25-04-2022,Barre au front derriere la tête,12,25.0,00:00:00
25-04-2022,Curl barre,12,30.0,00:00:00
25-04-2022,Barre au front derriere la tête,12,25.0,00:00:00
25-04-2022,Barre au front derriere la tête,12,25.0,00:00:00
25-04-2022,Curl barre,12,30.0,00:00:00
25-04-2022,Curl barre,12,30.0,00:00:00